hello
siva garu
march 25th 2025
